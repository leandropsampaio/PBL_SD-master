// Nios.v

// Generated using ACDS version 13.1 162 at 2018.11.06.09:36:31

`timescale 1 ps / 1 ps
module Nios (
		input  wire       clk_clk,                               //                            clk.clk
		output wire       led_external_connection_export,        //        led_external_connection.export
		input  wire       pushbuton1_external_connection_export, // pushbuton1_external_connection.export
		output wire       led2_external_connection_export,       //       led2_external_connection.export
		output wire       led3_external_connection_export,       //       led3_external_connection.export
		output wire       led4_external_connection_export,       //       led4_external_connection.export
		output wire       led5_external_connection_export,       //       led5_external_connection.export
		input  wire       pushbuton2_external_connection_export, // pushbuton2_external_connection.export
		input  wire       pushbuton3_external_connection_export, // pushbuton3_external_connection.export
		input  wire       pushbuton4_external_connection_export, // pushbuton4_external_connection.export
		output wire       lcd_rs,                                //                            lcd.rs
		output wire       lcd_rw,                                //                               .rw
		output wire       lcd_en,                                //                               .en
		output wire [7:0] lcd_db,                                //                               .db
		input  wire       uart_rxd,                              //                           uart.rxd
		output wire       uart_txd                               //                               .txd
	);

	wire         nios_jtag_debug_module_reset_reset;                                      // Nios:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios_custom_instruction_master_result;                                   // Nios_custom_instruction_master_translator:ci_slave_result -> Nios:E_ci_result
	wire   [4:0] nios_custom_instruction_master_b;                                        // Nios:D_ci_b -> Nios_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_c;                                        // Nios:D_ci_c -> Nios_custom_instruction_master_translator:ci_slave_c
	wire         nios_custom_instruction_master_done;                                     // Nios_custom_instruction_master_translator:ci_slave_multi_done -> Nios:E_ci_multi_done
	wire         nios_custom_instruction_master_clk_en;                                   // Nios:E_ci_multi_clk_en -> Nios_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] nios_custom_instruction_master_a;                                        // Nios:D_ci_a -> Nios_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_n;                                        // Nios:D_ci_n -> Nios_custom_instruction_master_translator:ci_slave_n
	wire         nios_custom_instruction_master_writerc;                                  // Nios:D_ci_writerc -> Nios_custom_instruction_master_translator:ci_slave_writerc
	wire         nios_custom_instruction_master_clk;                                      // Nios:E_ci_multi_clock -> Nios_custom_instruction_master_translator:ci_slave_multi_clk
	wire         nios_custom_instruction_master_reset_req;                                // Nios:E_ci_multi_reset_req -> Nios_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios_custom_instruction_master_start;                                    // Nios:E_ci_multi_start -> Nios_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] nios_custom_instruction_master_dataa;                                    // Nios:E_ci_dataa -> Nios_custom_instruction_master_translator:ci_slave_dataa
	wire         nios_custom_instruction_master_readra;                                   // Nios:D_ci_readra -> Nios_custom_instruction_master_translator:ci_slave_readra
	wire         nios_custom_instruction_master_reset;                                    // Nios:E_ci_multi_reset -> Nios_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] nios_custom_instruction_master_datab;                                    // Nios:E_ci_datab -> Nios_custom_instruction_master_translator:ci_slave_datab
	wire         nios_custom_instruction_master_readrb;                                   // Nios:D_ci_readrb -> Nios_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_result;        // Nios_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_b;             // Nios_custom_instruction_master_translator:multi_ci_master_b -> Nios_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_c;             // Nios_custom_instruction_master_translator:multi_ci_master_c -> Nios_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_a;             // Nios_custom_instruction_master_translator:multi_ci_master_a -> Nios_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk_en;        // Nios_custom_instruction_master_translator:multi_ci_master_clken -> Nios_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         nios_custom_instruction_master_translator_multi_ci_master_done;          // Nios_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios_custom_instruction_master_translator_multi_ci_master_n;             // Nios_custom_instruction_master_translator:multi_ci_master_n -> Nios_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         nios_custom_instruction_master_translator_multi_ci_master_writerc;       // Nios_custom_instruction_master_translator:multi_ci_master_writerc -> Nios_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk;           // Nios_custom_instruction_master_translator:multi_ci_master_clk -> Nios_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset_req;     // Nios_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios_custom_instruction_master_translator_multi_ci_master_start;         // Nios_custom_instruction_master_translator:multi_ci_master_start -> Nios_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_dataa;         // Nios_custom_instruction_master_translator:multi_ci_master_dataa -> Nios_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios_custom_instruction_master_translator_multi_ci_master_readra;        // Nios_custom_instruction_master_translator:multi_ci_master_readra -> Nios_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset;         // Nios_custom_instruction_master_translator:multi_ci_master_reset -> Nios_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_datab;         // Nios_custom_instruction_master_translator:multi_ci_master_datab -> Nios_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         nios_custom_instruction_master_translator_multi_ci_master_readrb;        // Nios_custom_instruction_master_translator:multi_ci_master_readrb -> Nios_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_result;         // Nios_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_b;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_c;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_done;           // Nios_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_a;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master0_n;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // Nios_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // Nios_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk;            // Nios_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // Nios_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_start;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readra;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_datab;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // Nios_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_result; // LCD_0:result -> Nios_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_start;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_start -> LCD_0:start
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> LCD_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_done;   // LCD_0:done -> Nios_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // Nios_custom_instruction_master_multi_slave_translator0:ci_master_clken -> LCD_0:clk_en
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_reset -> LCD_0:reset
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_datab -> LCD_0:datab
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // Nios_custom_instruction_master_multi_slave_translator0:ci_master_clk -> LCD_0:clk
	wire         nios_instruction_master_waitrequest;                                     // mm_interconnect_0:Nios_instruction_master_waitrequest -> Nios:i_waitrequest
	wire  [16:0] nios_instruction_master_address;                                         // Nios:i_address -> mm_interconnect_0:Nios_instruction_master_address
	wire         nios_instruction_master_read;                                            // Nios:i_read -> mm_interconnect_0:Nios_instruction_master_read
	wire  [31:0] nios_instruction_master_readdata;                                        // mm_interconnect_0:Nios_instruction_master_readdata -> Nios:i_readdata
	wire   [1:0] mm_interconnect_0_pushbuton4_s1_address;                                 // mm_interconnect_0:pushbuton4_s1_address -> pushbuton4:address
	wire  [31:0] mm_interconnect_0_pushbuton4_s1_readdata;                                // pushbuton4:readdata -> mm_interconnect_0:pushbuton4_s1_readdata
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                   // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire  [12:0] mm_interconnect_0_memory_s1_address;                                     // mm_interconnect_0:memory_s1_address -> memory:address
	wire         mm_interconnect_0_memory_s1_chipselect;                                  // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire         mm_interconnect_0_memory_s1_clken;                                       // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_memory_s1_write;                                       // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                    // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                  // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire  [15:0] mm_interconnect_0_uart_1_s1_writedata;                                   // mm_interconnect_0:UART_1_s1_writedata -> UART_1:writedata
	wire   [2:0] mm_interconnect_0_uart_1_s1_address;                                     // mm_interconnect_0:UART_1_s1_address -> UART_1:address
	wire         mm_interconnect_0_uart_1_s1_chipselect;                                  // mm_interconnect_0:UART_1_s1_chipselect -> UART_1:chipselect
	wire         mm_interconnect_0_uart_1_s1_write;                                       // mm_interconnect_0:UART_1_s1_write -> UART_1:write_n
	wire         mm_interconnect_0_uart_1_s1_read;                                        // mm_interconnect_0:UART_1_s1_read -> UART_1:read_n
	wire  [15:0] mm_interconnect_0_uart_1_s1_readdata;                                    // UART_1:readdata -> mm_interconnect_0:UART_1_s1_readdata
	wire         mm_interconnect_0_uart_1_s1_begintransfer;                               // mm_interconnect_0:UART_1_s1_begintransfer -> UART_1:begintransfer
	wire         mm_interconnect_0_nios_jtag_debug_module_waitrequest;                    // Nios:jtag_debug_module_waitrequest -> mm_interconnect_0:Nios_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_writedata;                      // mm_interconnect_0:Nios_jtag_debug_module_writedata -> Nios:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios_jtag_debug_module_address;                        // mm_interconnect_0:Nios_jtag_debug_module_address -> Nios:jtag_debug_module_address
	wire         mm_interconnect_0_nios_jtag_debug_module_write;                          // mm_interconnect_0:Nios_jtag_debug_module_write -> Nios:jtag_debug_module_write
	wire         mm_interconnect_0_nios_jtag_debug_module_read;                           // mm_interconnect_0:Nios_jtag_debug_module_read -> Nios:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_readdata;                       // Nios:jtag_debug_module_readdata -> mm_interconnect_0:Nios_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios_jtag_debug_module_debugaccess;                    // mm_interconnect_0:Nios_jtag_debug_module_debugaccess -> Nios:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios_jtag_debug_module_byteenable;                     // mm_interconnect_0:Nios_jtag_debug_module_byteenable -> Nios:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_led4_s1_writedata;                                     // mm_interconnect_0:led4_s1_writedata -> led4:writedata
	wire   [1:0] mm_interconnect_0_led4_s1_address;                                       // mm_interconnect_0:led4_s1_address -> led4:address
	wire         mm_interconnect_0_led4_s1_chipselect;                                    // mm_interconnect_0:led4_s1_chipselect -> led4:chipselect
	wire         mm_interconnect_0_led4_s1_write;                                         // mm_interconnect_0:led4_s1_write -> led4:write_n
	wire  [31:0] mm_interconnect_0_led4_s1_readdata;                                      // led4:readdata -> mm_interconnect_0:led4_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuton2_s1_address;                                 // mm_interconnect_0:pushbuton2_s1_address -> pushbuton2:address
	wire  [31:0] mm_interconnect_0_pushbuton2_s1_readdata;                                // pushbuton2:readdata -> mm_interconnect_0:pushbuton2_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuton1_s1_address;                                 // mm_interconnect_0:pushbuton1_s1_address -> pushbuton1:address
	wire  [31:0] mm_interconnect_0_pushbuton1_s1_readdata;                                // pushbuton1:readdata -> mm_interconnect_0:pushbuton1_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuton3_s1_address;                                 // mm_interconnect_0:pushbuton3_s1_address -> pushbuton3:address
	wire  [31:0] mm_interconnect_0_pushbuton3_s1_readdata;                                // pushbuton3:readdata -> mm_interconnect_0:pushbuton3_s1_readdata
	wire  [31:0] mm_interconnect_0_led3_s1_writedata;                                     // mm_interconnect_0:led3_s1_writedata -> led3:writedata
	wire   [1:0] mm_interconnect_0_led3_s1_address;                                       // mm_interconnect_0:led3_s1_address -> led3:address
	wire         mm_interconnect_0_led3_s1_chipselect;                                    // mm_interconnect_0:led3_s1_chipselect -> led3:chipselect
	wire         mm_interconnect_0_led3_s1_write;                                         // mm_interconnect_0:led3_s1_write -> led3:write_n
	wire  [31:0] mm_interconnect_0_led3_s1_readdata;                                      // led3:readdata -> mm_interconnect_0:led3_s1_readdata
	wire  [31:0] mm_interconnect_0_led2_s1_writedata;                                     // mm_interconnect_0:led2_s1_writedata -> led2:writedata
	wire   [1:0] mm_interconnect_0_led2_s1_address;                                       // mm_interconnect_0:led2_s1_address -> led2:address
	wire         mm_interconnect_0_led2_s1_chipselect;                                    // mm_interconnect_0:led2_s1_chipselect -> led2:chipselect
	wire         mm_interconnect_0_led2_s1_write;                                         // mm_interconnect_0:led2_s1_write -> led2:write_n
	wire  [31:0] mm_interconnect_0_led2_s1_readdata;                                      // led2:readdata -> mm_interconnect_0:led2_s1_readdata
	wire  [31:0] mm_interconnect_0_led5_s1_writedata;                                     // mm_interconnect_0:led5_s1_writedata -> led5:writedata
	wire   [1:0] mm_interconnect_0_led5_s1_address;                                       // mm_interconnect_0:led5_s1_address -> led5:address
	wire         mm_interconnect_0_led5_s1_chipselect;                                    // mm_interconnect_0:led5_s1_chipselect -> led5:chipselect
	wire         mm_interconnect_0_led5_s1_write;                                         // mm_interconnect_0:led5_s1_write -> led5:write_n
	wire  [31:0] mm_interconnect_0_led5_s1_readdata;                                      // led5:readdata -> mm_interconnect_0:led5_s1_readdata
	wire  [31:0] mm_interconnect_0_led1_s1_writedata;                                     // mm_interconnect_0:led1_s1_writedata -> led1:writedata
	wire   [1:0] mm_interconnect_0_led1_s1_address;                                       // mm_interconnect_0:led1_s1_address -> led1:address
	wire         mm_interconnect_0_led1_s1_chipselect;                                    // mm_interconnect_0:led1_s1_chipselect -> led1:chipselect
	wire         mm_interconnect_0_led1_s1_write;                                         // mm_interconnect_0:led1_s1_write -> led1:write_n
	wire  [31:0] mm_interconnect_0_led1_s1_readdata;                                      // led1:readdata -> mm_interconnect_0:led1_s1_readdata
	wire         nios_data_master_waitrequest;                                            // mm_interconnect_0:Nios_data_master_waitrequest -> Nios:d_waitrequest
	wire  [31:0] nios_data_master_writedata;                                              // Nios:d_writedata -> mm_interconnect_0:Nios_data_master_writedata
	wire  [16:0] nios_data_master_address;                                                // Nios:d_address -> mm_interconnect_0:Nios_data_master_address
	wire         nios_data_master_write;                                                  // Nios:d_write -> mm_interconnect_0:Nios_data_master_write
	wire         nios_data_master_read;                                                   // Nios:d_read -> mm_interconnect_0:Nios_data_master_read
	wire  [31:0] nios_data_master_readdata;                                               // mm_interconnect_0:Nios_data_master_readdata -> Nios:d_readdata
	wire         nios_data_master_debugaccess;                                            // Nios:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:Nios_data_master_debugaccess
	wire   [3:0] nios_data_master_byteenable;                                             // Nios:d_byteenable -> mm_interconnect_0:Nios_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;             // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                 // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         irq_mapper_receiver0_irq;                                                // UART_1:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_d_irq_irq;                                                          // irq_mapper:sender_irq -> Nios:d_irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [Nios:reset_n, UART_1:reset_n, irq_mapper:reset, led1:reset_n, led2:reset_n, led3:reset_n, led4:reset_n, led5:reset_n, memory:reset, mm_interconnect_0:Nios_reset_n_reset_bridge_in_reset_reset, pushbuton1:reset_n, pushbuton2:reset_n, pushbuton3:reset_n, pushbuton4:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [Nios:reset_req, memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset]

	Nios_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	Nios_Nios nios (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (nios_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios_data_master_read),                                //                          .read
		.d_readdata                            (nios_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios_data_master_write),                               //                          .write
		.d_writedata                           (nios_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios_instruction_master_read),                         //                          .read
		.i_readdata                            (nios_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (nios_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (nios_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (nios_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (nios_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (nios_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (nios_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (nios_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (nios_custom_instruction_master_reset_req)              //                          .reset_req
	);

	Nios_led1 led1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led1_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)        // external_connection.export
	);

	Nios_pushbuton1 pushbuton1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pushbuton1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuton1_s1_readdata), //                    .readdata
		.in_port  (pushbuton1_external_connection_export)     // external_connection.export
	);

	Nios_led1 led2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led2_s1_readdata),   //                    .readdata
		.out_port   (led2_external_connection_export)       // external_connection.export
	);

	Nios_led1 led3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led3_s1_readdata),   //                    .readdata
		.out_port   (led3_external_connection_export)       // external_connection.export
	);

	Nios_led1 led4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led4_s1_readdata),   //                    .readdata
		.out_port   (led4_external_connection_export)       // external_connection.export
	);

	Nios_led1 led5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_led5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led5_s1_readdata),   //                    .readdata
		.out_port   (led5_external_connection_export)       // external_connection.export
	);

	Nios_pushbuton1 pushbuton2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pushbuton2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuton2_s1_readdata), //                    .readdata
		.in_port  (pushbuton2_external_connection_export)     // external_connection.export
	);

	Nios_pushbuton1 pushbuton3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pushbuton3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuton3_s1_readdata), //                    .readdata
		.in_port  (pushbuton3_external_connection_export)     // external_connection.export
	);

	Nios_pushbuton1 pushbuton4 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pushbuton4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuton4_s1_readdata), //                    .readdata
		.in_port  (pushbuton4_external_connection_export)     // external_connection.export
	);

	lcd_driver lcd_0 (
		.datab  (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  // nios_custom_instruction_slave.datab
		.clk    (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                              .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.reset  (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.dataa  (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //                              .dataa
		.done   (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.result (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.rs     (lcd_rs),                                                                  //                   conduit_end.export
		.rw     (lcd_rw),                                                                  //                              .export
		.en     (lcd_en),                                                                  //                              .export
		.db     (lcd_db)                                                                   //                              .export
	);

	Nios_UART_1 uart_1 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_1_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_1_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_1_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_1_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_1_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_1_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_1_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_rxd),                                  // external_connection.export
		.txd           (uart_txd),                                  //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	Nios_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                    //                .ipending
		.ci_slave_estatus          (),                                                                    //                .estatus
		.ci_slave_multi_clk        (nios_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                    //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                    //                .datab
		.comb_ci_master_result     (),                                                                    //                .result
		.comb_ci_master_n          (),                                                                    //                .n
		.comb_ci_master_readra     (),                                                                    //                .readra
		.comb_ci_master_readrb     (),                                                                    //                .readrb
		.comb_ci_master_writerc    (),                                                                    //                .writerc
		.comb_ci_master_a          (),                                                                    //                .a
		.comb_ci_master_b          (),                                                                    //                .b
		.comb_ci_master_c          (),                                                                    //                .c
		.comb_ci_master_ipending   (),                                                                    //                .ipending
		.comb_ci_master_estatus    (),                                                                    //                .estatus
		.multi_ci_master_clk       (nios_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_result     (),                                                                    //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                         //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                             //     (terminated)
	);

	Nios_Nios_custom_instruction_master_multi_xconnect nios_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (nios_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	Nios_mm_interconnect_0 mm_interconnect_0 (
		.Clk_clk_clk                                   (clk_clk),                                                     //                                 Clk_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // jtag_uart_0_reset_reset_bridge_in_reset.reset
		.Nios_reset_n_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                              //      Nios_reset_n_reset_bridge_in_reset.reset
		.Nios_data_master_address                      (nios_data_master_address),                                    //                        Nios_data_master.address
		.Nios_data_master_waitrequest                  (nios_data_master_waitrequest),                                //                                        .waitrequest
		.Nios_data_master_byteenable                   (nios_data_master_byteenable),                                 //                                        .byteenable
		.Nios_data_master_read                         (nios_data_master_read),                                       //                                        .read
		.Nios_data_master_readdata                     (nios_data_master_readdata),                                   //                                        .readdata
		.Nios_data_master_write                        (nios_data_master_write),                                      //                                        .write
		.Nios_data_master_writedata                    (nios_data_master_writedata),                                  //                                        .writedata
		.Nios_data_master_debugaccess                  (nios_data_master_debugaccess),                                //                                        .debugaccess
		.Nios_instruction_master_address               (nios_instruction_master_address),                             //                 Nios_instruction_master.address
		.Nios_instruction_master_waitrequest           (nios_instruction_master_waitrequest),                         //                                        .waitrequest
		.Nios_instruction_master_read                  (nios_instruction_master_read),                                //                                        .read
		.Nios_instruction_master_readdata              (nios_instruction_master_readdata),                            //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.led1_s1_address                               (mm_interconnect_0_led1_s1_address),                           //                                 led1_s1.address
		.led1_s1_write                                 (mm_interconnect_0_led1_s1_write),                             //                                        .write
		.led1_s1_readdata                              (mm_interconnect_0_led1_s1_readdata),                          //                                        .readdata
		.led1_s1_writedata                             (mm_interconnect_0_led1_s1_writedata),                         //                                        .writedata
		.led1_s1_chipselect                            (mm_interconnect_0_led1_s1_chipselect),                        //                                        .chipselect
		.led2_s1_address                               (mm_interconnect_0_led2_s1_address),                           //                                 led2_s1.address
		.led2_s1_write                                 (mm_interconnect_0_led2_s1_write),                             //                                        .write
		.led2_s1_readdata                              (mm_interconnect_0_led2_s1_readdata),                          //                                        .readdata
		.led2_s1_writedata                             (mm_interconnect_0_led2_s1_writedata),                         //                                        .writedata
		.led2_s1_chipselect                            (mm_interconnect_0_led2_s1_chipselect),                        //                                        .chipselect
		.led3_s1_address                               (mm_interconnect_0_led3_s1_address),                           //                                 led3_s1.address
		.led3_s1_write                                 (mm_interconnect_0_led3_s1_write),                             //                                        .write
		.led3_s1_readdata                              (mm_interconnect_0_led3_s1_readdata),                          //                                        .readdata
		.led3_s1_writedata                             (mm_interconnect_0_led3_s1_writedata),                         //                                        .writedata
		.led3_s1_chipselect                            (mm_interconnect_0_led3_s1_chipselect),                        //                                        .chipselect
		.led4_s1_address                               (mm_interconnect_0_led4_s1_address),                           //                                 led4_s1.address
		.led4_s1_write                                 (mm_interconnect_0_led4_s1_write),                             //                                        .write
		.led4_s1_readdata                              (mm_interconnect_0_led4_s1_readdata),                          //                                        .readdata
		.led4_s1_writedata                             (mm_interconnect_0_led4_s1_writedata),                         //                                        .writedata
		.led4_s1_chipselect                            (mm_interconnect_0_led4_s1_chipselect),                        //                                        .chipselect
		.led5_s1_address                               (mm_interconnect_0_led5_s1_address),                           //                                 led5_s1.address
		.led5_s1_write                                 (mm_interconnect_0_led5_s1_write),                             //                                        .write
		.led5_s1_readdata                              (mm_interconnect_0_led5_s1_readdata),                          //                                        .readdata
		.led5_s1_writedata                             (mm_interconnect_0_led5_s1_writedata),                         //                                        .writedata
		.led5_s1_chipselect                            (mm_interconnect_0_led5_s1_chipselect),                        //                                        .chipselect
		.memory_s1_address                             (mm_interconnect_0_memory_s1_address),                         //                               memory_s1.address
		.memory_s1_write                               (mm_interconnect_0_memory_s1_write),                           //                                        .write
		.memory_s1_readdata                            (mm_interconnect_0_memory_s1_readdata),                        //                                        .readdata
		.memory_s1_writedata                           (mm_interconnect_0_memory_s1_writedata),                       //                                        .writedata
		.memory_s1_byteenable                          (mm_interconnect_0_memory_s1_byteenable),                      //                                        .byteenable
		.memory_s1_chipselect                          (mm_interconnect_0_memory_s1_chipselect),                      //                                        .chipselect
		.memory_s1_clken                               (mm_interconnect_0_memory_s1_clken),                           //                                        .clken
		.Nios_jtag_debug_module_address                (mm_interconnect_0_nios_jtag_debug_module_address),            //                  Nios_jtag_debug_module.address
		.Nios_jtag_debug_module_write                  (mm_interconnect_0_nios_jtag_debug_module_write),              //                                        .write
		.Nios_jtag_debug_module_read                   (mm_interconnect_0_nios_jtag_debug_module_read),               //                                        .read
		.Nios_jtag_debug_module_readdata               (mm_interconnect_0_nios_jtag_debug_module_readdata),           //                                        .readdata
		.Nios_jtag_debug_module_writedata              (mm_interconnect_0_nios_jtag_debug_module_writedata),          //                                        .writedata
		.Nios_jtag_debug_module_byteenable             (mm_interconnect_0_nios_jtag_debug_module_byteenable),         //                                        .byteenable
		.Nios_jtag_debug_module_waitrequest            (mm_interconnect_0_nios_jtag_debug_module_waitrequest),        //                                        .waitrequest
		.Nios_jtag_debug_module_debugaccess            (mm_interconnect_0_nios_jtag_debug_module_debugaccess),        //                                        .debugaccess
		.pushbuton1_s1_address                         (mm_interconnect_0_pushbuton1_s1_address),                     //                           pushbuton1_s1.address
		.pushbuton1_s1_readdata                        (mm_interconnect_0_pushbuton1_s1_readdata),                    //                                        .readdata
		.pushbuton2_s1_address                         (mm_interconnect_0_pushbuton2_s1_address),                     //                           pushbuton2_s1.address
		.pushbuton2_s1_readdata                        (mm_interconnect_0_pushbuton2_s1_readdata),                    //                                        .readdata
		.pushbuton3_s1_address                         (mm_interconnect_0_pushbuton3_s1_address),                     //                           pushbuton3_s1.address
		.pushbuton3_s1_readdata                        (mm_interconnect_0_pushbuton3_s1_readdata),                    //                                        .readdata
		.pushbuton4_s1_address                         (mm_interconnect_0_pushbuton4_s1_address),                     //                           pushbuton4_s1.address
		.pushbuton4_s1_readdata                        (mm_interconnect_0_pushbuton4_s1_readdata),                    //                                        .readdata
		.UART_1_s1_address                             (mm_interconnect_0_uart_1_s1_address),                         //                               UART_1_s1.address
		.UART_1_s1_write                               (mm_interconnect_0_uart_1_s1_write),                           //                                        .write
		.UART_1_s1_read                                (mm_interconnect_0_uart_1_s1_read),                            //                                        .read
		.UART_1_s1_readdata                            (mm_interconnect_0_uart_1_s1_readdata),                        //                                        .readdata
		.UART_1_s1_writedata                           (mm_interconnect_0_uart_1_s1_writedata),                       //                                        .writedata
		.UART_1_s1_begintransfer                       (mm_interconnect_0_uart_1_s1_begintransfer),                   //                                        .begintransfer
		.UART_1_s1_chipselect                          (mm_interconnect_0_uart_1_s1_chipselect)                       //                                        .chipselect
	);

	Nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (nios_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
